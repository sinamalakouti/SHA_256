library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Adder is
  Port (
  i , clk : in std_logic;
  o :out std_logic
         );
end Adder;
architecture Behavioral of q5 is 
end Behavioral;
