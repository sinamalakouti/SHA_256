library ieee;
use ieee.std_logic_1164.all;
use work.types.all;

package constants is

  constant pre_a : std_logic_vector(31 downto 0);
	constant pre_b : std_logic_vector(31 downto 0);
	constant pre_c : std_logic_vector(31 downto 0);
	constant pre_d : std_logic_vector(31 downto 0);
	constant pre_e : std_logic_vector(31 downto 0);
	constant pre_f : std_logic_vector(31 downto 0);
	constant pre_g : std_logic_vector(31 downto 0);
	constant pre_h : std_logic_vector(31 downto 0);

  constant k_values : K;

end package;

package body constants is
  constant pre_a : std_logic_vector(31 downto 0) := "01101010000010011110011001100111"; -- 6a09e667
	constant pre_b : std_logic_vector(31 downto 0) := "10111011011001111010111010000101"; -- bb67ae85
	constant pre_c : std_logic_vector(31 downto 0) := "00111100011011101111001101110010"; -- 3c6ef372
	constant pre_d : std_logic_vector(31 downto 0) := "10100101010011111111010100111010"; -- a54ff53a
	constant pre_e : std_logic_vector(31 downto 0) := "01010001000011100101001001111111"; -- 510e527f
	constant pre_f : std_logic_vector(31 downto 0) := "10011011000001010110100010001100"; -- 9b05688c
	constant pre_g : std_logic_vector(31 downto 0) := "00011111100000111101100110101011"; -- 1f83d9ab
	constant pre_h : std_logic_vector(31 downto 0) := "01011011111000001100110100011001"; -- 5be0cd19

  constant k_values : K := (
      "01000010100010100010111110011000", --428a2f98
      "01110001001101110100010010010001", --71374491
      "10110101110000001111101111001111", --b5c0fbcf
      "11101001101101011101101110100101", --e9b5dba5
      "00111001010101101100001001011011", --3956c25b
      "01011001111100010001000111110001", --59f111f1
      "10010010001111111000001010100100", --923f82a4
      "10101011000111000101111011010101", --ab1c5ed5
      "11011000000001111010101010011000", --d807aa98
      "00010010100000110101101100000001", --12835b01
      "00100100001100011000010110111110", --243185be
      "01010101000011000111110111000011", --550c7dc3
      "01110010101111100101110101110100", --72be5d74
      "10000000110111101011000111111110", --80deb1fe
      "10011011110111000000011010100111", --9bdc06a7
      "11000001100110111111000101110100", --c19bf174
      "11100100100110110110100111000001", --e49b69c1
      "11101111101111100100011110000110", --efbe4786
      "00001111110000011001110111000110", --0fc19dc6
      "00100100000011001010000111001100", --240ca1cc
      "00101101111010010010110001101111", --2de92c6f
      "01001010011101001000010010101010", --4a7484aa
      "01011100101100001010100111011100", --5cb0a9dc
      "01110110111110011000100011011010", --76f988da
      "10011000001111100101000101010010", --983e5152
      "10101000001100011100011001101101", --a831c66d
      "10110000000000110010011111001000", --b00327c8
      "10111111010110010111111111000111", --bf597fc7
      "11000110111000000000101111110011", --c6e00bf3
      "11010101101001111001000101000111", --d5a79147
      "00000110110010100110001101010001", --06ca6351
      "00010100001010010010100101100111", --14292967
      "00100111101101110000101010000101", --27b70a85
      "00101110000110110010000100111000", --2e1b2138
      "01001101001011000110110111111100", --4d2c6dfc
      "01010011001110000000110100010011", --53380d13
      "01100101000010100111001101010100", --650a7354
      "01110110011010100000101010111011", --766a0abb
      "10000001110000101100100100101110", --81c2c92e
      "10010010011100100010110010000101", --92722c85
      "10100010101111111110100010100001", --a2bfe8a1
      "10101000000110100110011001001011", --a81a664b
      "11000010010010111000101101110000", --c24b8b70
      "11000111011011000101000110100011", --c76c51a3
      "11010001100100101110100000011001", --d192e819
      "11010110100110010000011000100100", --d6990624
      "11110100000011100011010110000101", --f40e3585
      "00010000011010101010000001110000", --106aa070
      "00011001101001001100000100010110", --19a4c116
      "00011110001101110110110000001000", --1e376c08
      "00100111010010000111011101001100", --2748774c
      "00110100101100001011110010110101", --34b0bcb5
      "00111001000111000000110010110011", --391c0cb3
      "01001110110110001010101001001010", --4ed8aa4a
      "01011011100111001100101001001111", --5b9cca4f
      "01101000001011100110111111110011", --682e6ff3
      "01110100100011111000001011101110", --748f82ee
      "01111000101001010110001101101111", --78a5636f
      "10000100110010000111100000010100", --84c87814
      "10001100110001110000001000001000", --8cc70208
      "10010000101111101111111111111010", --90befffa
      "10100100010100000110110011101011", --a4506ceb
      "10111110111110011010001111110111", --bef9a3f7
      "11000110011100010111100011110010"  --c67178f2
		);
end package body;
